package shared_package;
	bit test_finished;
	integer Correct_counts = 0 ;
    integer Error_counts   = 0 ;
endpackage 